module module1 #(parameter DATA_WIDTH=1, DATA2 =3)(
    input [DATA_WIDTH-1:0] data_in,
    output [DATA2:0] data_out,
    output data_out_2,
    input  clk,
    input  rst,
);

endmodule;
