module module1 #(parameter DATA_WIDTH=1, DATA2 =3)(
    input [DATA_WIDTH-1:0] data_in, data_in_num_2, 
    output [DATA2:0] data_out, 
    input  clk,
    input  rst
);

endmodule;
