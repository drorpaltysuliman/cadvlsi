module module2(
    input [DATA_W2-1:0] data_in,
    output [2:0] data_out,
    output data_en,
    input  clk, clk_en,
    input  rst
);

endmodule;
