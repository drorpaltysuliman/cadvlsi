module block_c();

module1 instance3();
module1 instance5();
module2 instance4();

endmodule
