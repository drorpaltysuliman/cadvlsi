//-----------------------------------------------------
// Design Name : uart 
// File Name   : uart.v
// Function    : Simple UART
// Coder       : Deepak Kumar Tala
//-----------------------------------------------------
module uart (
// Port declarations
input        reset          ,
input        txclk          ,
input        ld_tx_data     ,
input  [7:0] tx_data        ,
input        tx_enable      );

//instance a 
// ggg sksks (

// AUTO_TEMPLATE check2(

//.bla(bla),
//.kjlds(uuduu));

// AUTO_TEMPLATE inst2c(
/*.input5(.*kkk));*/


check1 check2 (
    .input1(wire1),
    .input2  (wire2) ,
    .input3  (wire3),
    .input4  (wire4)   
);

inst2c #(.param1(uuud),.param2(mmsms[rr + 11pp])) check4 (
    .input1(wire1[5:4]),
    .input2  (wire2[PARAM2-1:0]) ,
    .input3  (wire3),
    .input4  (wire4)   
);

endmodule



